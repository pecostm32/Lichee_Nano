// Verilog netlist created by TD v5.0.28716
// Wed Apr  6 10:53:49 2022

`timescale 1ns / 1ps
module SIN_ROM  // sin_table.v(14)
  (
  addra,
  addrb,
  clka,
  clkb,
  rsta,
  rstb,
  doa,
  dob
  );

  input [11:0] addra;  // sin_table.v(21)
  input [11:0] addrb;  // sin_table.v(22)
  input clka;  // sin_table.v(23)
  input clkb;  // sin_table.v(24)
  input rsta;  // sin_table.v(25)
  input rstb;  // sin_table.v(26)
  output [13:0] doa;  // sin_table.v(18)
  output [13:0] dob;  // sin_table.v(19)


  // address_offset=0;data_offset=0;depth=4096;width=2;num_section=1;width_per_section=2;section_size=14;working_depth=4096;working_width=2;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h762DD887621D887721DC87722DC8B722DC8B722DD8B762DD8B762DD8B762DD88),
    .INIT_01(256'hDC8B7621DC8B762DD887722DC8B7621DC87722DD8B7621D887721DC8B722DD8B),
    .INIT_02(256'h77221DC8877221DC8877221DC8B7622DD8877221DC8B7621DC8B7621DC8B7621),
    .INIT_03(256'h8777222DDD88B776221DD88877622DDD88B77221DD88B77221DD88B7722DDC88),
    .INIT_04(256'h88888777762222DDDDC888877772222DDDC888B7772221DDD8887776221DDD88),
    .INIT_05(256'hB77777777777777777762222222222DDDDDDDDC8888888777777622222DDDDDC),
    .INIT_06(256'h778888888DDDDDDDD22222222227777777777777777778888888888888888888),
    .INIT_07(256'h22377488DDD222777888DDD22237778889DDDE222377748888DDDDD222223777),
    .INIT_08(256'hD22748DE23789DE27789DE23788DD227788DD227788DD2237488DD22377889DD),
    .INIT_09(256'h49E278D2349E278DE378D2348D2348D2378DE3789D2748DE2789D23789D23789),
    .INIT_0A(256'h49279E38D349E78D349E78D249E349278D278D249E349E349E348D278D278DE3),
    .INIT_0B(256'h4934E39E4934E39E4924D38E39E79E49249249249249249249249E79E78E34D3),
    .INIT_0C(256'h939393934E4E4E393938E4E493934E4E3938E4D3934E4938E4D39E4D39E4938E),
    .INIT_0D(256'h4E4E9393E4E4F9393A4E4E4F93939393E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E3),
    .INIT_0E(256'h90E90E90E90E53E53A4394E90E53A4F90E5394E93A4E93A4E93A4E5390E4F939),
    .INIT_0F(256'h0FE943E940FA50FA50FA50FA43E943E50FA43E90FA43E50E94FA43A53E50E90E),
    .INIT_10(256'hFEA95400FEA95403FAA5403FA9500FEA540FE9503FA540FA940FA940FA943EA5),
    .INIT_11(256'h555555540000000000003FFFFFFAAAAA955540003FFFAAA955400FFFAA95500F),
    .INIT_12(256'h00556ABFC00556AAFFC00555AAABFFF00015555AAAAAFFFFFFC0000000000001),
    .INIT_13(256'hF05AF05AF056BC16AF056BC05ABC05ABC056BF015ABF015ABF0156AFF0156ABF),
    .INIT_14(256'h6C1BC6B16C1AC5BC6B06B06B06B06B06BC5BC1AC16F05BC1AF05BC16B05AF05A),
    .INIT_15(256'hB1B1B1B1B1B1B1B1B1B1B16C6C6C6B1B1BC6C6F1B1AC6F1B06C5B1AC6B1AC5B1),
    .INIT_16(256'h1861B6DB2CB1C61B6CB186DB1C6DB1C6CB1B6C6DB1B6C6C71B1B2C6C6C6DB1B1),
    .INIT_17(256'h872DCB62D8721CB61CB61CB61CB61CB2D871CB6D871CB2DB6D861861C71C71C6),
    .INIT_18(256'h2DDDC888777222DDC8877622DD887722DD8B762DD8B721D8B721D8B72DC8721C),
    .INIT_19(256'h27778889DDDE2222777774888888889DDDDDDDDDDDDDDC88888888B777776222),
    .INIT_1A(256'hD278D2349D2789E2789E2749D23789D23789DE27789DE237489DE2277889DDE2),
    .INIT_1B(256'hE4D38E7924934D38E38E38E38E38E38D349249E38D349E38D278E349E349E348),
    .INIT_1C(256'h4E93939393939393939393939393938E4E4E793934E4E3938E4D3924E3924E39),
    .INIT_1D(256'h3E50E90E90E90E90E93E53A4394E93E4390E4390E4393E4E9390E4E539394E4E),
    .INIT_1E(256'hFFA9503FA540FE9503EA50FE940FA503E943E943E943E943E50FA43E90F943A5),
    .INIT_1F(256'hFFFFFFFFFFFFFFAAAAAA555540003FFFAAA555003FFAA95403FEA95403FAA540),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x14_sub_000000_000 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n8,open_n9,open_n10,1'b0,open_n11,open_n12,1'b0,open_n13,open_n14}),
    .dib({open_n15,open_n16,open_n17,1'b0,open_n18,open_n19,1'b0,open_n20,open_n21}),
    .rsta(rsta),
    .rstb(rstb),
    .doa({open_n26,open_n27,open_n28,open_n29,open_n30,open_n31,open_n32,doa[1:0]}),
    .dob({open_n33,open_n34,open_n35,open_n36,open_n37,open_n38,open_n39,dob[1:0]}));
  // address_offset=0;data_offset=2;depth=4096;width=2;num_section=1;width_per_section=2;section_size=14;working_depth=4096;working_width=2;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hD2749E378D2349D2789E378D2349D2789E378D2349D2789E378D2349D2789E34),
    .INIT_01(256'hE348D2789E378D2349E278DE348D2789E378D2349D278DE348D2749E278DE348),
    .INIT_02(256'hD278DE349D278DE349D278DE348D2789E348D2789E378D2749E278D2349D278D),
    .INIT_03(256'h48D278DE349E278D2789E349D278DE349E278D2749E378D2789E348D2789E349),
    .INIT_04(256'h49E348D278D2789E349E349D278D2789E349E378D278D2349E348D278D2349E3),
    .INIT_05(256'hD278D278D278D278D278D278D278D2349E349E349E349E278D278D278DE349E3),
    .INIT_06(256'h8D349E349E349E349278D278D278D278D278D278D278D349E349E349E349E349),
    .INIT_07(256'h8D278E349E38D278D349E34D278D279E349E34D278D279E349E349E78D278D27),
    .INIT_08(256'h4D279E34D279E34D279E34D279E34D278E349278D349E78D249E34D278D349E3),
    .INIT_09(256'h49E78E38D349279E38D34D249E78E34D279E38D349279E34D249E78D349278E3),
    .INIT_0A(256'h34D249249249E79E79E38E38E34D34D249279E79E38E34D349249E78E38D3492),
    .INIT_0B(256'h9E79E79E4924924934D34D34D34D34E38E38E38E38E38E38E38E34D34D34D34D),
    .INIT_0C(256'h924D38E79E4934D38E79E4934D38E39E7924934D38E39E79E4924934D34E38E3),
    .INIT_0D(256'h4934E7924E39E4D38E4934E3924D38E7934E39E4934E39E4934E39E4934E39E7),
    .INIT_0E(256'h4E3934E4939E4D3924E7934E4938E4939E4D39E4D39E4D39E4D39E4D39E4938E),
    .INIT_0F(256'hE393924E4E3939E4E493934E4D3938E4E3938E4E3938E4E3934E4D3924E4939E),
    .INIT_10(256'h4E4E4E4E39393938E4E4E4D393939E4E4E49393924E4E493939E4E4E393924E4),
    .INIT_11(256'h4E4E4E4E4E4E4E4E4E4E7939393939393939393924E4E4E4E4E4E3939393939E),
    .INIT_12(256'h4E4E4E4E5393939393A4E4E4E4E4E4E93939393939393939390E4E4E4E4E4E4E),
    .INIT_13(256'h3E4E439394E4E539394E4E539390E4E4F939394E4E4E939393E4E4E4E9393939),
    .INIT_14(256'h3A4E5394E5390E4F93E4E9394E4393E4E5390E4F9394E4F9394E4F9394E4E939),
    .INIT_15(256'hE93E4394E93E4394E93E4390E53A4E93E4F90E4394E5394E93A4E93A4E93A4E9),
    .INIT_16(256'h90E93E53E53E53E43A43A4F94F90E90E53E43A4F94E90E53E4394F90E53A4394),
    .INIT_17(256'hF94FA43E50E94F943A43E53E90E94F94FA43A43A53E53E53E50E90E90E90E90E),
    .INIT_18(256'h3A50FA50E943E90FA50E943E50FA43E90FA43E90FA43E90F943E50E94FA53E90),
    .INIT_19(256'hE943FA50FA503E943E943FA50FA50FA50FA50FA50FA50FA50FA50F943E943E94),
    .INIT_1A(256'h03EA543FA543FA543FA543FA543EA503E950FA943FA503E950FA543E950FA503),
    .INIT_1B(256'h00FEA5403FA9503FA9503FA9503FA9503FA950FEA540FA9503EA540FA950FEA5),
    .INIT_1C(256'hFAA95403FEA95403FEA95403FEA9540FFAA5403FEA5503FEA5503FEA5403FA95),
    .INIT_1D(256'h3FFFAAA555000FFFAA9554003FFAA955400FFEAA55403FFAA95500FFEA95500F),
    .INIT_1E(256'hAAAAAA955555000003FFFFAAAAA555540003FFFEAAA95554000FFFEAAA555400),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAAAAAAAAAA955555555400000003FFFFFF),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x14_sub_000000_002 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n48,open_n49,open_n50,1'b0,open_n51,open_n52,1'b0,open_n53,open_n54}),
    .dib({open_n55,open_n56,open_n57,1'b0,open_n58,open_n59,1'b0,open_n60,open_n61}),
    .rsta(rsta),
    .rstb(rstb),
    .doa({open_n66,open_n67,open_n68,open_n69,open_n70,open_n71,open_n72,doa[3:2]}),
    .dob({open_n73,open_n74,open_n75,open_n76,open_n77,open_n78,open_n79,dob[3:2]}));
  // address_offset=0;data_offset=4;depth=4096;width=2;num_section=1;width_per_section=2;section_size=14;working_depth=4096;working_width=2;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h543FA543FA940FA940FA940FE950FE950FE9503EA503EA503EA543FA543FA540),
    .INIT_01(256'hFEA503EA503EA543FA543FA540FA940FA940FE950FE950FEA503EA503EA503FA),
    .INIT_02(256'h543FA540FA940FA950FE950FEA503EA503FA543FA543FA940FA940FE950FE950),
    .INIT_03(256'hFA543FA540FA940FE950FEA503EA503FA543FA940FA940FE950FEA503EA503FA),
    .INIT_04(256'h0FA950FE9503EA503FA540FA940FE950FEA503EA543FA940FA950FE9503EA503),
    .INIT_05(256'h03EA543FA940FE9503EA543FA940FE950FEA503FA540FA940FE9503EA503FA54),
    .INIT_06(256'h0FEA503FA540FA9503EA543FA940FE9503EA543FA940FEA503FA540FA950FEA5),
    .INIT_07(256'hFA940FEA503FA940FEA503FA940FE9503FA540FE9503EA540FA950FEA543FA94),
    .INIT_08(256'h503EA540FE9503FA940FEA543FA9503EA540FE9503FA540FEA503FA940FEA503),
    .INIT_09(256'hA503FA9503FA940FEA540FEA503FA9503EA540FEA543FA9503FA540FEA543FA9),
    .INIT_0A(256'h9503FA9503FA540FEA540FEA540FEA540FE9503FA9503FA9503FA540FEA540FE),
    .INIT_0B(256'h0FEA540FFA9503FA9503FA9503FA9503FA9503FA9503FA9503FA9503FA9503FA),
    .INIT_0C(256'h540FEA540FFA9503FA9500FEA540FEA5403FA9503FA9503FAA540FEA540FEA54),
    .INIT_0D(256'h503FA9540FEA5503FAA540FEA9503FA9540FEA5503FA9500FEA540FFA9503FA9),
    .INIT_0E(256'hFA9540FFA9500FEA9503FEA5503FAA540FFA9500FEA5503FAA540FFA9500FEA5),
    .INIT_0F(256'hFEA9540FFA9540FFAA5403FAA5403FAA5403FAA5403FAA5403FAA5403FAA540F),
    .INIT_10(256'hA5500FFA95403FEA5500FFA95403FAA5500FEA9540FFAA5403FAA5503FEA9500),
    .INIT_11(256'hFAA5500FFAA5500FFAA5403FEA95403FEA95403FEA5500FFAA5503FEA95403FA),
    .INIT_12(256'hA5500FFAA95403FEA95500FFAA5500FFEA95403FEA95403FEAA5500FFAA5500F),
    .INIT_13(256'hEAA55403FFAA55403FFAA55403FFAA55003FEAA5500FFEA95400FFAA55403FEA),
    .INIT_14(256'h955003FFAA95500FFEAA55400FFEA955003FFAA55400FFAA95500FFEAA55003F),
    .INIT_15(256'hAA955400FFEAA955003FFEAA55400FFEAA555003FFAA955003FFAA955003FFAA),
    .INIT_16(256'h55003FFEAA9554003FFEAA555000FFFAA955400FFFAAA554003FFAAA554003FF),
    .INIT_17(256'h5550003FFFAAA5554003FFEAAA555000FFFEAA9554003FFEAAA555000FFFAAA5),
    .INIT_18(256'h3FFFAAAA5554000FFFFAAA95550003FFFAAA95550003FFFAAA9555000FFFEAAA),
    .INIT_19(256'hFFFEAAAA555540003FFFEAAAA55550000FFFFAAAA55550000FFFFAAA95554000),
    .INIT_1A(256'h5400003FFFFEAAAA95555400003FFFFEAAAA5555400003FFFFAAAA9555500003),
    .INIT_1B(256'h00FFFFFFEAAAAA9555554000003FFFFFEAAAAA555555000003FFFFFAAAAA5555),
    .INIT_1C(256'h00000003FFFFFFFEAAAAAAA9555555500000003FFFFFFEAAAAAA955555540000),
    .INIT_1D(256'hEAAAAAAAAAAAA5555555555540000000000FFFFFFFFFEAAAAAAAAA5555555550),
    .INIT_1E(256'hAAAAAAAAAAAAAAAAA9555555555555555554000000000000000FFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAAAAA),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x14_sub_000000_004 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n88,open_n89,open_n90,1'b0,open_n91,open_n92,1'b0,open_n93,open_n94}),
    .dib({open_n95,open_n96,open_n97,1'b0,open_n98,open_n99,1'b0,open_n100,open_n101}),
    .rsta(rsta),
    .rstb(rstb),
    .doa({open_n106,open_n107,open_n108,open_n109,open_n110,open_n111,open_n112,doa[5:4]}),
    .dob({open_n113,open_n114,open_n115,open_n116,open_n117,open_n118,open_n119,dob[5:4]}));
  // address_offset=0;data_offset=6;depth=4096;width=2;num_section=1;width_per_section=2;section_size=14;working_depth=4096;working_width=2;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h003FFFFEAAAAA5555500000FFFFFAAAAA55555400003FFFFEAAAA95555400000),
    .INIT_01(256'h000003FFFFEAAAA95555400000FFFFFAAAAA5555500000FFFFFEAAAA95555400),
    .INIT_02(256'h55400000FFFFFAAAAA55555000003FFFFEAAAA95555400000FFFFFAAAAA55555),
    .INIT_03(256'h5555400000FFFFFAAAAA55555400003FFFFEAAAAA5555500000FFFFFEAAAA955),
    .INIT_04(256'hA55555000003FFFFEAAAAA5555500000FFFFFEAAAA95555500000FFFFFEAAAA9),
    .INIT_05(256'hA95555400000FFFFFEAAAA95555500000FFFFFEAAAAA55555000003FFFFEAAAA),
    .INIT_06(256'hA55555400000FFFFFEAAAA955555000003FFFFEAAAAA55555400000FFFFFAAAA),
    .INIT_07(256'h55555000003FFFFFAAAAA955555000003FFFFFAAAAA95555500000FFFFFEAAAA),
    .INIT_08(256'h55400000FFFFFEAAAAA555554000003FFFFFAAAAA955555000003FFFFFAAAAA9),
    .INIT_09(256'h0003FFFFFEAAAAA555555000003FFFFFEAAAAA555554000003FFFFFAAAAA9555),
    .INIT_0A(256'hFFFEAAAAA955555000000FFFFFFAAAAAA555554000003FFFFFEAAAAA55555500),
    .INIT_0B(256'hA5555550000003FFFFFEAAAAA9555554000003FFFFFEAAAAA9555554000003FF),
    .INIT_0C(256'h000FFFFFFAAAAAA9555555000000FFFFFFEAAAAA9555554000000FFFFFFAAAAA),
    .INIT_0D(256'hAA95555550000003FFFFFFAAAAAA95555550000003FFFFFFAAAAAA5555554000),
    .INIT_0E(256'hFFFFFFAAAAAAA55555540000003FFFFFFAAAAAAA5555554000000FFFFFFFAAAA),
    .INIT_0F(256'h0000000FFFFFFFAAAAAAA955555540000003FFFFFFEAAAAAA95555554000000F),
    .INIT_10(256'h5555500000003FFFFFFFAAAAAAA955555550000000FFFFFFFEAAAAAA95555555),
    .INIT_11(256'h555555500000000FFFFFFFEAAAAAAA9555555540000000FFFFFFFEAAAAAAA955),
    .INIT_12(256'h55555000000003FFFFFFFFAAAAAAAA55555555400000003FFFFFFFFAAAAAAAA5),
    .INIT_13(256'h00000003FFFFFFFFEAAAAAAAA955555555400000000FFFFFFFFFAAAAAAAA9555),
    .INIT_14(256'hFFFFFEAAAAAAAAA55555555550000000003FFFFFFFFFAAAAAAAAA55555555540),
    .INIT_15(256'h5555555500000000003FFFFFFFFFFAAAAAAAAAA955555555540000000003FFFF),
    .INIT_16(256'hFFFFEAAAAAAAAAAA95555555555500000000000FFFFFFFFFFFEAAAAAAAAAA955),
    .INIT_17(256'h0000003FFFFFFFFFFFFEAAAAAAAAAAAA5555555555554000000000000FFFFFFF),
    .INIT_18(256'h400000000000000FFFFFFFFFFFFFFEAAAAAAAAAAAAA955555555555550000000),
    .INIT_19(256'h00000000000000003FFFFFFFFFFFFFFFFAAAAAAAAAAAAAAAA555555555555555),
    .INIT_1A(256'h0000003FFFFFFFFFFFFFFFFFFFEAAAAAAAAAAAAAAAAAA9555555555555555554),
    .INIT_1B(256'hFFAAAAAAAAAAAAAAAAAAAAAAAA95555555555555555555555400000000000000),
    .INIT_1C(256'h555555540000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA55555555555555555555555555555),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAAAAAAAAAAA),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x14_sub_000000_006 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n128,open_n129,open_n130,1'b0,open_n131,open_n132,1'b0,open_n133,open_n134}),
    .dib({open_n135,open_n136,open_n137,1'b0,open_n138,open_n139,1'b0,open_n140,open_n141}),
    .rsta(rsta),
    .rstb(rstb),
    .doa({open_n146,open_n147,open_n148,open_n149,open_n150,open_n151,open_n152,doa[7:6]}),
    .dob({open_n153,open_n154,open_n155,open_n156,open_n157,open_n158,open_n159,dob[7:6]}));
  // address_offset=0;data_offset=8;depth=4096;width=2;num_section=1;width_per_section=2;section_size=14;working_depth=4096;working_width=2;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFEAAAAAAAAAAAAAAAAAAAA55555555555555555555400000000000000000000),
    .INIT_01(256'hAAAAA95555555555555555555500000000000000000000FFFFFFFFFFFFFFFFFF),
    .INIT_02(256'h55555555000000000000000000003FFFFFFFFFFFFFFFFFFFFAAAAAAAAAAAAAAA),
    .INIT_03(256'h0000000000FFFFFFFFFFFFFFFFFFFFEAAAAAAAAAAAAAAAAAAAA5555555555555),
    .INIT_04(256'hFFFFFFFFFFFEAAAAAAAAAAAAAAAAAAAA55555555555555555555500000000000),
    .INIT_05(256'hAAAAAAAAAAAA5555555555555555555550000000000000000000003FFFFFFFFF),
    .INIT_06(256'h5555555555550000000000000000000003FFFFFFFFFFFFFFFFFFFFFAAAAAAAAA),
    .INIT_07(256'h00000000003FFFFFFFFFFFFFFFFFFFFFEAAAAAAAAAAAAAAAAAAAAA5555555555),
    .INIT_08(256'hFFFFFFFFAAAAAAAAAAAAAAAAAAAAAA9555555555555555555555400000000000),
    .INIT_09(256'hAAA95555555555555555555555400000000000000000000003FFFFFFFFFFFFFF),
    .INIT_0A(256'h000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFEAAAAAAAAAAAAAAAAAAA),
    .INIT_0B(256'hFFFFFFFFFFFFFEAAAAAAAAAAAAAAAAAAAAAAA955555555555555555555555400),
    .INIT_0C(256'hAAA55555555555555555555555550000000000000000000000000FFFFFFFFFFF),
    .INIT_0D(256'h0000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFEAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_0E(256'hAAAAAAAAAAAAAAAAAAAAAAAAAA95555555555555555555555555500000000000),
    .INIT_0F(256'h555555500000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFA),
    .INIT_10(256'hFFFFFFFFFFFFEAAAAAAAAAAAAAAAAAAAAAAAAAAAAA5555555555555555555555),
    .INIT_11(256'h5555555555555550000000000000000000000000000000FFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFEAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA955555555555555555),
    .INIT_13(256'h5555555400000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA955555555555555555555555555555),
    .INIT_15(256'h0000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAAA),
    .INIT_16(256'h5555555555555555555555555555555555555550000000000000000000000000),
    .INIT_17(256'hFFFFFFEAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA5555555),
    .INIT_18(256'h000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h5555555555555555400000000000000000000000000000000000000000000000),
    .INIT_1A(256'hAAAAAA9555555555555555555555555555555555555555555555555555555555),
    .INIT_1B(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x14_sub_000000_008 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n168,open_n169,open_n170,1'b0,open_n171,open_n172,1'b0,open_n173,open_n174}),
    .dib({open_n175,open_n176,open_n177,1'b0,open_n178,open_n179,1'b0,open_n180,open_n181}),
    .rsta(rsta),
    .rstb(rstb),
    .doa({open_n186,open_n187,open_n188,open_n189,open_n190,open_n191,open_n192,doa[9:8]}),
    .dob({open_n193,open_n194,open_n195,open_n196,open_n197,open_n198,open_n199,dob[9:8]}));
  // address_offset=0;data_offset=10;depth=4096;width=2;num_section=1;width_per_section=2;section_size=14;working_depth=4096;working_width=2;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h5555555555555555555555555555555555555555555555000000000000000000),
    .INIT_02(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAA955555555555555555555555555555555555),
    .INIT_03(256'hFFFFFFFFFFAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000003FFFFFFFFF),
    .INIT_06(256'h5555555555555555555555555555555554000000000000000000000000000000),
    .INIT_07(256'hAAAAAAAAAA955555555555555555555555555555555555555555555555555555),
    .INIT_08(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAAAAAAAAAAAAA),
    .INIT_0A(256'h000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h5555555555555555555555555555555555555555555555555555500000000000),
    .INIT_0D(256'hAAAAAAAAAAAAAAA9555555555555555555555555555555555555555555555555),
    .INIT_0E(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h0000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFF),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h5555555555555555555555555555555555555555555000000000000000000000),
    .INIT_14(256'h5555555555555555555555555555555555555555555555555555555555555555),
    .INIT_15(256'hAAAAAAAAAAAAAAAAAA9555555555555555555555555555555555555555555555),
    .INIT_16(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_17(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_18(256'hFFFFFFFFFFFFFFFAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x14_sub_000000_010 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n208,open_n209,open_n210,1'b0,open_n211,open_n212,1'b0,open_n213,open_n214}),
    .dib({open_n215,open_n216,open_n217,1'b0,open_n218,open_n219,1'b0,open_n220,open_n221}),
    .rsta(rsta),
    .rstb(rstb),
    .doa({open_n226,open_n227,open_n228,open_n229,open_n230,open_n231,open_n232,doa[11:10]}),
    .dob({open_n233,open_n234,open_n235,open_n236,open_n237,open_n238,open_n239,dob[11:10]}));
  // address_offset=0;data_offset=12;depth=4096;width=2;num_section=1;width_per_section=2;section_size=14;working_depth=4096;working_width=2;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  AL_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h5555555555555555555555555555555555555555555555555555554000000000),
    .INIT_06(256'h5555555555555555555555555555555555555555555555555555555555555555),
    .INIT_07(256'h5555555555555555555555555555555555555555555555555555555555555555),
    .INIT_08(256'h5555555555555555555555555555555555555555555555555555555555555555),
    .INIT_09(256'h5555555555555555555555555555555555555555555555555555555555555555),
    .INIT_0A(256'hAAAAAAAAAAAAAAAAAAAAA5555555555555555555555555555555555555555555),
    .INIT_0B(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_0C(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_0D(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_0E(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_0F(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_10(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAAAAAAAAAAAAAAAA),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_4096x14_sub_000000_012 (
    .addra({addra,1'b1}),
    .addrb({addrb,1'b1}),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n248,open_n249,open_n250,1'b0,open_n251,open_n252,1'b0,open_n253,open_n254}),
    .dib({open_n255,open_n256,open_n257,1'b0,open_n258,open_n259,1'b0,open_n260,open_n261}),
    .rsta(rsta),
    .rstb(rstb),
    .doa({open_n266,open_n267,open_n268,open_n269,open_n270,open_n271,open_n272,doa[13:12]}),
    .dob({open_n273,open_n274,open_n275,open_n276,open_n277,open_n278,open_n279,dob[13:12]}));

endmodule 

